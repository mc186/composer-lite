module adder (input reg [31:0] a,
              input reg [31:0] b,
              output reg [31:0] c);

  assign c= a + b;
endmodule

